typedef enum bit[1:0] {
    FIXED,
    INCR,
    WRAP
  } burst_type_t;
  
  `define DATA_WIDTH 32
  `define ADDR_WIDTH 16
